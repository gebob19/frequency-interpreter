module main (
	// Inputs
	CLOCK_50,
	SW,
	KEY,
	AUD_ADCDAT,

	// Bidirectionals
	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,
	I2C_SDAT,

	// Outputs
	AUD_XCK,
	AUD_DACDAT,
	I2C_SCLK,
	VGA_CLK,   						//	VGA Clock
	VGA_HS,							//	VGA H_SYNC
	VGA_VS,							//	VGA V_SYNC
	VGA_BLANK_N,					//	VGA BLANK
	VGA_SYNC_N,						//	VGA SYNC
	VGA_R,   						//	VGA Red[9:0]
	VGA_G,	 						//	VGA Green[9:0]
	VGA_B,
	HEX0,
	HEX1,
	HEX2,
	HEX3,
	HEX4,
	HEX5,
	HEX6,
	HEX7,
	LEDR,
	LEDG
);
	// Inputs
	input				CLOCK_50;
    input [9:0] SW;
    input [3:0] KEY;
	input				AUD_ADCDAT;

	// Bidirectionals
	inout				AUD_BCLK;
	inout				AUD_ADCLRCK;
	inout				AUD_DACLRCK;
	inout				I2C_SDAT;

	// Outputs
	output				AUD_XCK;
	output				AUD_DACDAT;
	output				I2C_SCLK;
	output 				VGA_CLK;   		//	VGA Clock
	output 				VGA_HS;			//	VGA H_SYNC
	output 				VGA_VS;			//	VGA V_SYNC
	output 				VGA_BLANK_N;	//	VGA BLANK
	output 				VGA_SYNC_N;		//	VGA SYNC
	output [9:0] VGA_R;   				//	VGA Red[9:0]
	output [9:0] VGA_G;	 				//	VGA Green[9:0]
	output [9:0] VGA_B;   				//	VGA Blue[9:0]

    output [17:0] LEDR;
    output [7:0] LEDG;
	output [6:0] HEX0;
	output [6:0] HEX1;
	output [6:0] HEX2;
	output [6:0] HEX3;
	output [6:0] HEX4;
	output [6:0] HEX5;
	output [6:0] HEX6;
	output [6:0] HEX7;

	// Internal Wires
	wire				audio_in_available;
	wire		[31:0]	left_channel_audio_in;
	wire		[31:0]	right_channel_audio_in;
	wire				read_audio_in;
	wire				audio_out_allowed;
	wire		[31:0]	left_channel_audio_out;
	wire		[31:0]	right_channel_audio_out;
	wire				write_audio_out;
	wire        [18:0]  delay;
	wire                tick;
	wire                reset;
	wire        [3:0]   frequency;
	wire [19199:0] image;
	wire [2:0] color_background;
	wire [2:0] color_foreground;

	// Internal Registers
	reg [18:0] delay_cnt;
	reg snd;
    reg [31:0] buff;
	reg [19199:0] current_image;
	reg [2:0] color_background_reg;
	reg [2:0] color_foreground_reg;

	/*****************************************************************************
	*                             Sequential Logic                              *
	*****************************************************************************/

	assign frequency = SW[3:0];
	assign delay = {frequency, 15'd3000};
	assign image = current_image;
	assign color_background = color_background_reg;
	assign color_foreground = color_foreground_reg;

	always @(posedge CLOCK_50)
	begin
		if(delay_cnt == delay) begin
			delay_cnt <= 0;
			snd <= !snd;
		end else delay_cnt <= delay_cnt + 1;
	end

	wire [27:0] sample_rate = 28'b10111110101111000001111111;

	ratedivider_28bit rateOne (
		.clock(CLOCK_50),
		.d(sample_rate),
		.enable(tick)
	);

	/*****************************************************************************
	*                            Combinational Logic                            *
	*****************************************************************************/

	assign resetn = KEY[0];

	wire [31:0] sound = (SW == 0) ? 0 : snd ? 32'd10000000 : -32'd10000000;

	assign read_audio_in			= audio_out_allowed;
	assign write_audio_out			= audio_out_allowed;
	assign left_channel_audio_out	= sound;
	assign right_channel_audio_out	= sound;

	always @(posedge tick) 
	begin
		buff <= sound;
	end

	/*****************************************************************************
	*                              Internal Modules                             *
	*****************************************************************************/

	Audio_Controller Audio_Controller (
		// Inputs
		.CLOCK_50						(CLOCK_50),
		.reset						(~resetn),

		.clear_audio_in_memory		(),
		.read_audio_in				(read_audio_in),
		
		.clear_audio_out_memory		(),
		.left_channel_audio_out		(left_channel_audio_out),
		.right_channel_audio_out	(right_channel_audio_out),
		.write_audio_out			(write_audio_out),

		.AUD_ADCDAT					(AUD_ADCDAT),

		// Bidirectionals
		.AUD_BCLK					(AUD_BCLK),
		.AUD_ADCLRCK				(AUD_ADCLRCK),
		.AUD_DACLRCK				(AUD_DACLRCK),


		// Outputs
		.audio_in_available			(audio_in_available),
		.left_channel_audio_in		(left_channel_audio_in),
		.right_channel_audio_in		(right_channel_audio_in),

		.audio_out_allowed			(audio_out_allowed),

		.AUD_XCK					(AUD_XCK),
		.AUD_DACDAT					(AUD_DACDAT),
	);

	/*****************************************************************************
	*                           Finite State Machine                             *
	*****************************************************************************/
    
    localparam STATE_LO3 = 4'b0000;
	localparam STATE_LO2 = 4'b0001;
	localparam STATE_LO1 = 4'b0011;
	localparam STATE_MEL = 4'b0010;
	localparam STATE_ME  = 4'b0110;
	localparam STATE_MEH = 4'b0100;
	localparam STATE_HI1 = 4'b1100;
	localparam STATE_HI2 = 4'b1000;
	localparam STATE_HI3 = 4'b1001;

	localparam INITIAL_STATE = STATE_ME;

	localparam TRANSITION_OFF = 2'b00;
	localparam TRANSITION_HI = 2'b01;
	localparam TRANSITION_ME = 2'b10;
	localparam TRANSITION_LO = 2'b11;

    reg [3:0] current_state, next_state;
    wire [1:0] transition;
	
	assign transition = (frequency + 4) / 5;

    always @(posedge tick)
    begin: state_table
        case (current_state)
            STATE_LO3:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_LO2;
						TRANSITION_ME: next_state <= STATE_LO2;
						TRANSITION_HI: next_state <= STATE_LO2;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b001;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000011111111111111111111100000000000000000000000000001111111111111111110000000000111111111111111000000000000000000001111111111111110000000000000000000000000000000001111111111111111111111000000000000000000000000000111111111111111111000000000011111111111111100000000000000000000111111111111111000000000000000000000000000000000001111111111111111111110000000000000000000000011111111111111111111100000000001111111111111111000000000000000000011111111111111110000000000000000000000000000000000111111111111111111111100000000000000000000111111111111111111111110000000000111111111111111110000000000000000001111111111111111000000000000000000001000000000000011111111111111111111111000000000000000000111111111111111111111111000000000011111111111111111000000000000000000011111111111111100000000000000000000011100000000000111111111111111111111111000000000000001111111111111111111111111000000000011111111111111111100000000000000000001111111111111110000000000000000000000000000000000000111111111111111111111111110000001111111111111111111111111111000000000001111111100011111110000000000000000000111111111111111100000000000000000010000110000000000001111111111111111111111111111111111111111111111111111111100000000000000111111000000111111100000000000000001111111111111111110000000000000000000000001001000110000011111111111111111111111111111111111111111111111111111110000000000000011111100000001111111011111111111111111111111111111111000000000000000000010000100100000000001111111111111111111111111111111111111111111111111111111000000000000001111110000000111111111111111111111111111111111111111100000000000000000000000000001110000000001111111111111111111111111111111111111111111111111111000000000000000111111000000011111111111111111111111111111111111111110000000000000000000000000000000010000000011111111111111111111111111111111111111111111110111001000000000000011111100000001111111111111111111111111111111111111111000000000000000000000000000000001000000000011111111111111111111111111111111111111111110010001101000000000001111110000000111111111111111111111111111111111111111100000000000000000000001000000000100000000001111111111111111111111111111111111111111111001001010000000000000111111000000011111111111111111111111111111111111000110000000000000000000000000000000100000000000011111111111111111111111111111111111111111110101100110000000000011111000000000111111111111111111111111111111111000011000000000000000000000001100000111000000000001111111111111111111111111111111111111111111001000010010000000001111100000000111111111111111111111111111111111000001100000000000000000000000111001111100000000000011111111111111111111111111111111111111111100000000001000000000111110000000011111111111111111111111111111111000100100000000000000000000000011111111110000000000000111111111111111111111111111111111111111000000000000100000000011100000000011111111111111111111111111111110000110100000000000000000000000001111111111000000000000111111111111111111111111111111111111110000001000000000000000011110000000000111111111111111111111111111110000111100000000000000000000000000111111111100000000000011111111111111111111111111111111111111000000000000000000001000000010000000111111111111111111111111111110000011100000000000000000000000000011111111110000000000001111111111111111111111111111111111111100000011000001000000100000000000000011111111111111111111111111110000001100000000000000000000000000000111111111000000000000011111111111111111111111111111111111110000001000000110000000000000010000011111111111111111111111110000000001100000000001000100000000000000001111111111000000000000001111111111111111111111111111111111000001111110110000000000000110000011111111111111111111111100000000111000000000010000000000000000000000011111111110000000000000011111111111111111111111111111111000000111111111000000000000110000111111111111111111111111100000000110000000000010000000000000000000000001111111111000000000000001111111111111111111111111111110000000011111111100000100000010001111111111111111111111111100000000110000000111100000110000000000000000000111111111100000000000000111111111111111111111111111111000000001111111110000010000010000111111111111111111111111111000000110000000110100000100000000000000000000011111111110000000000000111111111111111111111111111111000000000111111111000010000010001111111111111111111111111111100001110000000110000000000000000000000000000000111111111110000000000011111111111111111111111111111100000000011111111000011000011111111111111111111111111111111000111000000011110000000000000000000000000000000001111111111110000000001111111111111111111111111111110000001111111111100011100011111111111111111111111111111111101111000000111110000000100000000000000000000000000111111111111100000000011111111111111111111111111110000000111111111110001100001011111111111111111111111111111111110000000111111000000100000000000000000000000000011111111111110000000011111111111111111111111111111100000111111111111001110000101111111111111111111111111111111110000000011111100000110000000000000000000000000000111111111111100000011111111111111111111111111111111000011111111111000100000010111111111111111111111111111111100000000011111110000000000000000000000000000000000000111111111111000011111111111111111111111111111111100011111111111000010000010011111111111111111111111111111110000000111000000010000000000000000000000000000000000011111111111100001111111111111111111111111111111110001111111111000000000001001111111111111111111111111111111000000111000000100000000000000000000000000000000000000011111111111111111111111111111111111111111111111000111111111100000000000100011111111111111111111111111111100000011100000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100111111111100000100000010001111111111111111111111111111111000011100000100000000000000000000000000000000000000000111111111111111111111111111111111111111111111110111111111110000010000001000111111111111111111111111111111100001110000010000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000001000000100011111111111111111111111111111110001111000100000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000100000010001111111111111111111111111111110000111000010000000000000000000000000000000000000000000001111111111111111111111111111111101111111111111111111111000000010000001000111111111111111111111111111111000111000010000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000001000000110011111111111111111111111111111100011000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111100000000000000001001111111111111111111111111111110011100001000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000001000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111110000000000100000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000010000111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111101111111111100000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111110111111111110000000001111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111000011111111111111100000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111001111111111111110000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111100000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111011100111111000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000111110001011011111100000000000000000000000000000001111111111111111110001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111000000000111110000000000000000000000000000000011111111111111111100111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111110000011111000000000000000000000000000000000001111111111111111000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111100000000000000000000000000000000000000111110111111110001111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000001111011111111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000001101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110001111111100000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000111110000000000000000000000000000000000000000000011011100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100111110000000000000000000000000000000000000000000011011110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000001111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000001101111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000110111110111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011011111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end
            STATE_LO2:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_LO3;
						TRANSITION_ME: next_state <= STATE_LO1;
						TRANSITION_HI: next_state <= STATE_LO1;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b001;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000011111111111111111000000000000000000000000011111111111111000000000000000011111111111111100000000000000011111111111111111110000000000000000000000000000000000000000111111111111111000000000000000000000000001111111111111000000000000000001111111111111110000000000000000011111111111111111100000000000000000000000000000000000000011111111111111100000000000000000000000000111111111111110000000000000000111111111111111000000000000000000111111111111111111000000000000000000000000000000000000000111111111111111000000000000000000000000011111111111111000000000000000111111100111111100000000000000000011111111111111111110000000000000000000000000000000000000001111111111111100000000000000000000000011111111111111100000000000000011111100000011110000000000000000000111111111111111111000000000000000000000000000000000000000111111111111110000000000000000000000001111111111111100000000000000001111110000000111000000000000000000001111111111111111100000000000000000000000000000000000000011111111111111000000000000000000000000111111111111110000000000000000011110000000011100000000000000000001111111111111111110000000000000000000000000000000000000001111111111111110000000000000000000000111111111111100000000000000000011111000000001110000000000000000011111111111111100010000000000000000000000000000000000000000011111111111111000000000000000000000111111111111110000000000000000000111100000000111100000000000000001111111111111100011100000000000000000000000000000000000000001111111111111110000000000000000000011111111111111000000000000000000011110000000011110000000000000001111111111111000001110000000000000000000000000000000000000000111111111111111000000000000000000011111111111111100000000000000000001111000000000111000000000000001111111111111000000110000000000000000000000000000000000000000001111111111111110000000000000000011111111111111100000000000000000000111100000000011100000000000001111111111111000000111000000000000000000000000000000000000000000111111111111111110000000000000011111111111111110000000000000000000011110000000001111000000000011111111111111000000111000000000000000000000000000000000000000000001111111111111111000000000000011111111111111110000000000000000000001111000000000111100000000011111111111111000000011000000000000000000000000000000000000000000000111111111111111110000000000111111111111111111000000000000000000000111100000000011110000000011111111111111000000011000000000000000000000000000000000000000000000011111111111111111100000000111111111111111111100000000000000000000011110000000001111100000111111111111111000000001000000000000000000000000000000000000000000000000111111111111111111110011111111111111111111110000000000000000000001111000000000111110000111111111111111000000011000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111000000000000000000000111100000000011111111111111111111111100000011100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000011110000000001111111111111111111111100000001100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111100000000000000000000001111000000000111111011111111111111110000001100000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000111100000000111111101111111111111110000000100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000011110000000011111100011111111111111000000100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000001111000000001111111111111111111111100000110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000111100000001111111111111111111111100000110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000011110000001111111111111111111111100000011000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000001111000000111111111111111111111110000011000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000111100000111111111111111111111100000010000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000011110000111111111111111111111110000010000000000000000000000000000000000000000000000110000000000000111111111111111111111111111111111111000000000000000000000000001111110111111111111111111111110001111000000000000000000000000000000000000000000000011111000000000011111111111111111111111111111111111110000000000100000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000110000000000001111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111110000011111111111111100000000000000000000000001111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111000000011111111111110000000000000000000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000001100000000000001111111111111111111111111111111110000110000000000000000000011111111111111111111111111111111100000000000000000000000001111000000000000000000100000110000000000000001111111111111111111111111111110000000000000000000000000001111111111111111111111111111111100000000000000000000000011000000000000000000000011111111000000000000000111111111111111111111111111111000000000000000000000000000001111111111111111111111111111100000000000000000111011000000000000000000000000001111111110000000000000001111111111111111111111111111000000000000000000000000000000111111111111111111111111111110000000000000011110000000000000000000000000000000111111111000000000000000111111111111111111111111111100000000000001000000000000000111111111111111111111111111110000000000001111110000000000000000000000000000000001111111110000000000000111111111111111111111111111100000000000000100000000000000111111111111111111111111111111000000000001111110000000000000000000000000000000000111111111000000000000111111111111111111111111111111000000000000010000000000000111111111111111111111111111111110000000001111111000000000000000000000000000000000011111111110000000000011111111111111111111111111111100000011111111000001100000011111111111111111111111111111111000000011111110100000000000000000000000000000000000111111111000000000001111111111111111111111111111100000001111111100000100000001111111111111111111111111111111100000011110000000110000000000000000000000000000000011111111100000000000011111111111111111111111111110000000111111110000110000110111111111111111111111111111111110000001110000000000000000000000000000000000000000001111111111000000000001111111111111111111111111111100000011111111000110000011011111111111111111111111111111111000001110000000011000000000000000000000000000000000011111111111000000000111111111111111111111111111110000101111111000011000000101111111111111111111111111111111100000100000000110000000000000000000000000000000000000111111111111000000111111111111111111111111111111100111111111100001100000010011111111111111111111111111111110000110000001100000000000000000000000000000000000000001111111111100000111111111111111111111111111111110011111111100000110000000101111111111111111111111111111111000111000001000000000000000000000000000000000000000000011111111110000011111111111111111111111111111111011111111110000011000000010111111111111111111111111111111100111100000100000000000000000000000000000000000000000001111111111100001111111111111111111111111111111001111111111000001100000001011111111111111111111111111111100011110000000000000000000000000000000000000000000000000011111111111100111111111111111111111111111111101111111111000000110000001101111111111111111111111111111100011100000010000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110111111111000000011000000011111111111111111111111111111110001110000001000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111011111111100000001100000001111111111111111111111111111111101111100001100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111110000000111000000111111111111111111111111111111111111111000100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000011101001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000001111111111111111000111111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111101111111111111100000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100011111111111000000000000000000000000000000011111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111001111111110000000000000000000000000000000000011111111111111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000111111100000000000000000000000000000000000000111110111111100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000010111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111001111100000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111100111110000000000000000000000000000000000000000000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110010000001111000000000000000000000000000000000000000000000011011110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111001000000111100000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100011111110000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111110000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010000011111000000000000000000000000000000000000000000011011111001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111000000000000000000000000000000000000000000001101111101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000111111110111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011100000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000001111100000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end
            STATE_LO1:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_LO2;
						TRANSITION_ME: next_state <= STATE_MEL;
						TRANSITION_HI: next_state <= STATE_MEL;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b001;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000000000011111111110000000000000000000000000011111111111000000000000000000001111111111111100000000000000111111111111111000000000000000000000000000000000000000000000000001111111111100000000000000000000000001111111111100000000000000000000111111111111110000000000000011111111111111100000000000000000000000000000000000000000000000000111111111110000000000000000000000000111111111110000000000000000000011111111111111100000000000001111111111111111000000000000000000000000000000000000000000000000011111111111000000000000000000000000011111111111000000000000000000001111111111111110000000000000011111111111111100000000000000000000000000000000000000000000000011111111111100000000000000000000000001111111111100000000000000000000111111111111111000000000000001111111111111110000000000000000000000000000000000000000000000001111111111111000000000000000000000000111111111110000000000000000000001111111111111100000000000000011111111111111000000000000000000000000000000000000000000000000111111111111100000000000000000000000111111111111000000000000000000000111111100001110000000000000001111111111111100000000000000000000000000000000000000000000000001111111111110000000000000000000000111111111111100000000000000000000011111100000111000000000000000111111111111111000000000000000000000000000000000000000000000000111111111111100000000000000000000111111111111110000000000000000000000111110000001100000000000000011111111111001110000000000000000000000000000000000000000000000001111111111111000000000000000000011111111111111000000000000000000000011110000000110000000000000111111111111000011000000000000000000000000000000000000000000000000111111111111110000000000000000001111111111111000000000000000000000011110000000001000000000000011111111111000001100000000000000000000000000000000000000000000000011111111111111000000000000000001111111111111100000000000000000000000111100000001100000000000001111111111000000110000000000000000000000000000000000000000000000000111111111111100000000000000000111111111111100000000000000000000000011110000000110000000000001111111111000000111000000000000000000000000000000000000000000000000011111111111110000000000000000011111111111110000000000000000000000001110000000011000000000000111111111100000011000000000000000000000000000000000000000000000000001111111111111000000000000000001111111111111000000000000000000000000111000000000100000000000111111111100000001100000000000000000000000000000000000000000000000000111111111111100000000000000001111111111111000000000000000000000000111100000000110000000000111111111100000001110000000000000000000000000000000000000000000000000001111111111110000000000000000111111111111100000000000000000000000011110000000011000000000011111111100000000110000000000000000000000000000000000000000000000000000111111111111000000000000000011111111111110000000000000000000000001111000000001100000000011111111110000000111000000000000000000000000000000000000000000000000000011111111111110000000000000001111111111111000000000000000000000000011100000000110000000011111111110000000011100000000000000000000000000000000000000000000000000001111111111111000000000000000111111111111100000000000000000000000011110000000011000000001111111111000000011110000000000000000000000000000000000000000000000000000011111111111110000000000000111111111111110000000000000000000000001111000000001100000001111111111000000001110000000000000000000000000000000000000000000000000000001111111111111000000000000011111111111111000000000000000000000000111100000000111000000111111111100000001111000000000000000000000000000000000000000000000000000000111111111111110000000000011111111111111100000000000000000000000011110000000011100000111111111100000000111000000000000000000000000000000000000000000000000000000011111111111111100000000011111111111111100000000000000000000000001110000000001110000111111111110000000111000000000000000000000000000000000000000000000000000000001111111111111111100000111111111111111110000000000000000000000000111000000001111111111111111111100000111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000011110000000111111111111111111110000011100000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000011111111000011111111111111111111000011110000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111101110000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000111111111111110011111111111111111100000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000001111111111110001111111111111111100000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111101000000000000000000000000000010111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000001001111111111111111111111111110000000000000000000000000000000000000000000000000000001110000000000000000001111111111111111111111111100000000000000000000000000000000111111111111111111111111111100000000000111111111111110000000000000000000000000001111110000000000000000111111111111111111111111110000000000000000000000100000001111111111111111111111111111110000000001111111111000000000000000000000000000000000100111100000000000000111111111111111111111111111000000000000000000000010000011111111111111111111111111111111000000001111111100000000000000000000000000000000000001001111000000000000011111111111111111111111111110000000100000000000011000001111111111111111111111111111111100000001111001110000000000000000000000000000000000000000111000000000000001111111111111111111111111111100001110000000000001000000011111111111111111111111111111110000001110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000001111111111111111111111111111111000001000000000001100000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000011111111111111111111111111111100001100000000000000000000000000000000000000000000011000001110000000000011111111111111111111111111111100000000000000000000000000001111111111111111111111111111110001110000000000000000000000000000000000000000000000111111111100000000001111111111111111111111111111110000010000100000000000000000111111111111111111111111111110000110000000000000000000000000000000000000000000000001111111111000000000011111111111111111111111111111000001000010000000000000000111111111111111111111111111111000111000000000000000000000000000000000000000000000000011111111100000000000111111111111111111111111111100001111111000000000000000011111111111111111111111111111000111000000000000000000000000000000000000000000000000001111111111100000000011111111111111111111111111110000111111100000000000000001111111111111111111111111111100111000000000000000000000000000000000000000000000000000011111111111000000011111111111111111111111111111001111111110000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111110000001111111111111111111111111111100111111111000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111100001111111111111111111111111111110111111111000000000011001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111000111111111111111111111111111110011111111000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111111111100011111111111111111111111111111001111111100000000011111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111100111111111111111111111111111101111111100000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111110111111110000000000011111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111111111100111111111111111111111111111111110000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111001111111111111111111111111111110000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111110111111111011111011111011111111000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111101111111111111101111101111111100000000000000000001111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000011111111111110111111111111110101000111111100000000000000000000011111111111111110001111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111011100010111110000000000000000000000011111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111010111011111000000000000000000000000011111111110110000011111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100111100111000000000000000000000000000011111111011100001111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110111110111100000000000000000000000000000011101011111000100000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111011111111100000000000000000000000000000000010001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111101111110000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000111001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000011111000000000000000000000000000000000000000000000001111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111001111000000000000000000000000000000000000000000000000101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000001110000000000000000000000000000000000000000000011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001111000111000000000000000000000000000000000000000000001101111001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000001100000000000000000000000000000000000000000000110111101111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000110000000000000000000000000000000000000000000011100000011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000111000000000000000000000000000000000000000000001111000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100011111100000000000000000000000000000000000000000000011100000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111110000000000000000000000000000000000000000000001111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000011100000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000011100000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101100011110000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end 
            STATE_MEL:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_LO1;
						TRANSITION_ME: next_state <= STATE_MEH;
						TRANSITION_HI: next_state <= STATE_MEH;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b010;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000000000000011111111100000000000000000000011111111000000000000000000011111111110000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000001111111000000000000000000001111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000111111110000000000000000000111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000111111111000000000000000000011111111110000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111100000000000000000001111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000111111110000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111000000000000000000001111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111100000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000111111110000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111110000000000000000000001111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111000000000000000000000111111111110000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111100000000000000000000011111111111000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000111111110000000000000000000001111111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111000000000000000000000111111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111000000000000000000000011111111111000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111100000000000000000000000111111111100000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001111111110000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000111111110000000000000000000000001111111111100000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000011111111000000000000000000000000111111111110000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000011111111100000000000000000000000001111111111000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000001111111110000000000000000000000000111111111100000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000001111111110000000000000000000000000011111111111000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000111111111000000000000000000000000001111111111100000111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000111111111100000000000000000000000000111111111110000011111111101000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111110000000000000000000000000011111111111100001111111100100000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000011111111111000000000000000000000000001111111111110000111111111010000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000111111111111000000000000000000000000000111111111111000011111111101000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000011111111111100000000000000000000000000011111111111110011111111110100000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000011111111111110000000000000000000000000001111111111111001111111111010000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100001111111111111000000000000000000000000000111111111111100111111111101000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110001111111111111100000000000000000000000000001111111111111011111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000011111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000111000000111111111111111111111111111111000000000000000000000000000111111111111111111111111110010000000000000000000000000000000000000000000000000000000000000000011100000011111111111111111111111111111100000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011100000001111111111111111111111111111110000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001100000000111111111111111111111111111111000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001110011000111111111111111111111111111111000000000000000000000000000111111111111111111111111110011000000000000000000000000000000000000000000000000000000000000000110000000011111111111111111111111111111100000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000010001000001111111111111111111111111111110000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001000000000011111111111111111111111111111100000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000100000000001111111111111111111111111111110000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011110000000111111111111111111111111111111000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111100000011111111111111111111111111111000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111110000001111111111100001111111111111100000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111000000111111111100011001111111111100000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111100000001111111111101111111111111100000000000000000000001000001001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111000000111111111111111111111111100000000000000000000000100000100111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111100000011111111111111111111111111000000000000000000000010000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111110000001111111111111111111111111100000000000000000000001000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111000000111111111111111111111111110000000000000000000000100000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111100000111111111111111111111111111000000000000000000000010000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111110000011111111111111111111111111100000000000000000000001000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111000001111111111111111111111111100000000000000000000000100000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111110000111111111111111111111111111000000000000000000000010000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111000011111111111111111111111111100000000000000000000001000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111100001111111111111111111111111110000000000000000000000100000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111110000011111111111111111111111111000000000000000000000010000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111000001111111111111111111111111100000000000000000000001000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111100000111111111111111111111111110000000000000000000000100000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111110000011111111111111111111111111100000000000000000000010000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000111111000000111111111111111111111111110000000000000000000001000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000011111110000011111111111111111111111111000000000000000000000100000100111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000001111111000001111111111111111111111111100000000000000000000010000010011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011111110001111111111111111111111111110000000000000000000001000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000001111111000111111111111111111111111111000000000000000000000100000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111111111111100000000000000000000010000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111111111110000000000000000000000011011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111111111111000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000001111111111111111111111011111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111100011100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000111111100111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111110011110111111111111111111111111111111111100000000001111111111111111111101111111111111111111111111111111000000000000000000000000000000000000000000000000000111111000001011011111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111110000001000011111111111111111111111111111000000000000111111111111111111111111111111111111111110000100110000000000000000000000000000000000000000000000000000111011100000110001111111110101111111111111111100000000000001111111111111111111111111111111111100000000010000000000000000000000000000000000000000000000000000000011101101001111001111110011000111111111111111110000000000000001111111111111111111111111111111100000000001000010000000000000000000000000000000000000000000000000000100011000111111111111011100111111100001111111000000000000000001111111100000011111000000000000000000000100001000000000000000000000000000000000000000000000000000000011111011111111111111111110111100000111111100000000000000000001111010011000110000000000000000000000010000100000000000000000000000000000000000000000000000000000000111011111111111111111111011100000011111110000000000000000000000000011110000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000001111111000000000000000000000000011111100000000000000000000000000010000100000000000000000000000000000000000000000000000000000000001111111111111111100000000000000111111100000000000000000000000011111111000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111110000000000000000000000001111111100000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000111111110111110000000000000001111111000000000000000000000000111000011000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000011111011001111000000000000000111111100000000000000000000000000001100000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000001111111000111100000000000000011111100000000000000000000000000011111100000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000111111111111110000000000000001111110000000000000000000000000000011000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001111111001111000000000000000111110000000000000000000000000000001110000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000110011110011100000000000000011111000000000000000000000000010000000000000000000000000000000000001011000000000000000000000000000000000000000000000000000000000000011000000001110000000000000001111100000000000000000000000011001000010010000000000000000000000000101100000000000000000000000000000000000000000000000000000000000011100000001111100000000000000111110000000000000000000000001101111011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110011111110000000000000010011000000000000000000000000110111101111100000000000000000000000001000100000000000000000000000000000000000000000000000000000000000111111101101110000000000000001001100000000000000000000000001100000000010000000000000000000000000010010000000000000000000000000000000000000000000000000000000000011101100010111000000000000001100110000000000000000000000000111100000111000000000000000000000000001110000000000000000000000000000000000000000000000000000000000001111000000111100000000000010000001000000000000000000000000011111000111110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000111111111111100000000000010000000100000000000000000000000000111111111111000000000000000000000001000001000000000000000000000000000000000000000000000000000000000011111111111110000000000010010000010000000000000000000000000011111111111000000000000000000000000101000100000000000000000000000000000000000000000000000000000000000111111111110000000000000001000000000000000000000000000000000011111111100000000000000000000000011000001000000000000000000000000000000000000000000000000000000000001111111111000000000000000100000000000000000000000000000000000011111100000000000000000000000001100000100000000000000000000000000000000000000000000000000000000000111111111000000000000000001010010000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000010100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end 
            STATE_ME:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_MEL;
						TRANSITION_ME: next_state <= STATE_ME;
						TRANSITION_HI: next_state <= STATE_MEH;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b010;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000000000000000001111111111000000000000000000000111111110000000000000000000111111111110000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000011111111000000000000000000001111111111000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000001111111100000000000000000000111111111100000000000111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000001111111110000000000000000000011111111110000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000111111111000000000000000000001111111111000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000011111111100000000000000000000111111111100000000000111111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000001111111110000000000000000000001111111110000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000111111110000000000000000000000111111111100000000001111111111100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000011111111000000000000000000000011111111110000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000001111111100000000000000000000001111111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000001111111110000000000000000000000111111111100000000001111111111100000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111110000000000000000000000011111111111000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111000000000000000000000001111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000000000000000000111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000001111111110000000000000000000000011111111111000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111000000000000000000000000111111111100000000011111111111000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111000000000000000000000000011111101110000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000011111111100000000000000000000000001111111111100000000111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000001111111110000000000000000000000000111111111110000000111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000111111110000000000000000000000000011111111111000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000111111111000000000000000000000000001111111111100000001111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000011111111100000000000000000000000000111111111110000000111111111001000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000011111111110000000000000000000000000011111111111100000011111111100100000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000001111111111000000000000000000000000001111111111110000011111111110010000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000001111111111100000000000000000000000000111111111111000001111111111011000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000111111111110000000000000000000000000011111111111110000111111111100100000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000111111111111000000000000000000000000001111111111111000011111111110010000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000111111111111000000000000000000000000000111111111111100011111111111001000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000011111111111100000000000000000000000000011111111111110001111111111100100000000000000000000000000000000000000000000000000000000000000000000000011111111111110000011111111111110000000000000000000000000001111111111111100111111111110010000000000000000000000000000000000000000000000000000000000000000000000001111111111111100001111111111111000000000000000000000000000111111111111110111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000111111111111100000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000011111111111111111111111111000100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000011111111111111111111111111001100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000011111111111111111111111110001100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000001111111111111111111111111100110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111110001111111111111100000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111110001100111111111100000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111110111111111111110000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000011111111111111111111111111110000000000000011111000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000010000000000000010000001111111111111111111111111110000000000000111111111111101110000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000011111100000111111111111111111111111111000000000001111111111110001000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000011111111000111111111111111111111111111100000000001111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111000000010000000001111111111111111111111111111111111111110000000011100000001100000000000000000000000000000000000000111110000000000000111111111111111111111111111100000011000000000011111110000000011111111111111111111111000100111100000000000000000000000000000000000000000000000111111110000000000011111111111111111111111111110000001100000000001000000000000001111111111111111111111100011111100000011110001110000000000000000000000000000011111111111111000000001111111111111111111111111110000001111000000000100000000000111111111111111111111111110011111100000111000000000000000000000000000000000000000100110000111111000000111111111111111111111111111000001111100010000001000000111111111111111111111111111111111111000000110000000000000000000000000000000000000001000000000111111111000011111111111111111111111111100001111111110000000100000011111111111111111111111111111111111110000010000000000000000000000000000000000000000010000000011111111111001111111111111111111111111111011111110010000000000000011111111111111111111111111111111111111100010000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000110011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111001111111111111111111111111111100000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111100001101101011111111111111111100000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000001111111110000000110101011111111111111110000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111111000000011000101111111011111110000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000111111111110011100111110110001111110000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111100101110111111101001111111000000000000000000000000000011111111110000111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111110111111000000000000000000000000000000111111110000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000110111111111111111111111111011000000000000000000000000000000000011101011100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111100000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100011110000000000000000000000000000000000000000000000011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001110011100000000000000000000000000000000000000000001000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000100001110000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110110001111100000000000000000000000000000000000000000001001110011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111110000000000000000000000000000000000000000000110111101011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111000000000000000000000000000000000000000000011100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000011100000000000000000000000000000000000000000000111000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000011100000000000000000000000000000000000000000000011111000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end 
            STATE_MEH:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_MEL;
						TRANSITION_ME: next_state <= STATE_MEL;
						TRANSITION_HI: next_state <= STATE_HI1;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b010;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000000000000000000000000001111111110000000000000000000001111111000000000000000000111111111100000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111100000000000000000001111111110000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000111111111000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111100000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111100000000000000000001111111110000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000111111110000000000000000000111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111000000000000000000011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111100000000000000000001111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000000000000000111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111110000000000000000000011111111110000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111110000000000000000000001111111111000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001111111000000000000000000000111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111100000000000000000000011111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111110000000000000000000001111111111000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111000000000000000000000111111111100000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000011111111100000000000000000000011111111110000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001111111100000000000000000000001111100111000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000111111110000000000000000000000011111111100000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000111111110000000000000000000000001111111111000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000011111111000000000000000000000000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000011111111100000000000000000000000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000001111111110000000000000000000000001111111111000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000001111111111000000000000000000000000111111111110000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000111111111100000000000000000000000001111111111000001111111101000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000111111111100000000000000000000000000111111111100000111111110110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000011111111110000000000000000000000000011111111110000011111111011000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000111111111111000000000000000000000000001111111111100011111111101100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000011111111111100000000000000000000000000111111111110001111111110110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000011111111111110000000000000000000000000011111111111100111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100001111111111110000000000000000000000000001111111111110011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111100000000000000000000000000111111111111011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000001111111111111111111111111110000000100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000111111111111111111111111111000000011000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000111111111111111111111111111100000010100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000011111111111111111111111111100000101000100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000010000000000000000011111111111111111111111111111000000110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000001111000000000000001111111111111111111111111111100000100010000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000100100000000000000011111111111111111111111111110000100001000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000011000000000000000001111111111111111111111110011000000000100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100010000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000101000000000000000000011111111111111111111111111100000100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000001000010000000000000001111111111111111111111111110000010010000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100001000000000000000000000111111111111111111111111111100001011000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000001100000000000000000011111111111111111111111111110000100000000000000000000000000000000000000000000000000000000000000000000000011111111111000111111111111110000001111100000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000110011111111111000000111110000000000000000111111111111111111111111111000010001000000000000000000000000000000000000000000000000000000000000000000000011111111111011111111111111000000011111000000000000000011111111111111111111111111100001000100000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110100000011111100000000000000001111111111111111111111111110000100010000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000001111110000000000000000111111111111111111111111110000010001000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000111111000000000000000011111111111111111111111111100011000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000111111100000000000000001111111111111111111111111110001000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000011111100000000000000000111111111111111111111111111000100010000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000001111110000000000000000011111111111111111111111111100110001000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100001111111000000000000000001111111111111111111111111110011000100000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110000111111000000000000000000111111111111111111111111111001100100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100011111100000000000000000011111111111111111111111111101100010000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110001111110000000000000000001111111111111111111111111110110001000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111001111111000000000000000000111111111111111111111111111011000100000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100111111000000000000000000011111111111111111111111111111100010000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110111111100000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111011111110000000000000000000111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000011111111111111111111111111111100010000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000001111111111111111111111111111100001000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000111111111111111111111111111110001000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000011111111111111111111111111111000100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000001111111111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000001100111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111111111111110111111111111111111111111110000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111111111111110011100111011111111110111111000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000001111111111111111111111111000011011001111111111011111000000000111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000001111111111111111111111111100100111100101100010001111100000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111110111011111111111001001111100000000000111110001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111000001010111111111110011111111111100111110110000000000011111000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111000000000000011111111110111111111111111110001000000000000110100000000001101111111110000001111100000000000000000000000000000000000000000000000000000000001111111100000000000000011111111111111111111111111000000000000000100001000000000000000110111110000110000000000000000000000000000000000000000000000000000000000000111111110000000000000000000001111111111111111111100000000000000000000100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000011111111111111110000000000000000000100010000000000000000001111111000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111111111110000000000000000000010001000000000000000000111111110000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000011111110011111000000000000000000001000000000000000000000111000111000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000001111111101111100000000000000000000100001000000000000000011011001100000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000111111100111110000000000000000000000000100000000000000000111111000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000011111111111111000000000000000000000100010000000000000000011100100000000000000000000000000000000000000000000000000000000000000000111001000000000000000000000000001111111101111100000000000000000000010001000000000000000000111100000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000111001100001110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000011100100000111000000000000000000000010010000000000000000111000000010000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000001100110011111100000000000000000000001000000000000000000011100111001000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000111111111111110000000000000000000000000100000000000000011111111000100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000011111111111110000000000000000000000001111000000000000001000000110010000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000001111100000111000000000000000000000000111110000000000000111000000111000000000000000000000000000000000000000000000000000000000001000111000000000000000000000000000111110000111100000000000000000000000010111000000000000011111111111100000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000011111111111100000000000000000000000000000100000000000001111111111100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111111110000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000011111111110000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000111111111000000000000000000000000001100001100000000000001111110000000000000000000000000000000000000000000000000000000000001000010010000000000000000000000000000011111111000000000000000000000000000011110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000011100000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000010101110000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000010011100000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end 
            STATE_HI1:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_MEH;
						TRANSITION_ME: next_state <= STATE_MEH;
						TRANSITION_HI: next_state <= STATE_HI2;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b100;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000000000001111111111000000000000000000000011111111100000000000000000000000000000111111111111000000000000000011111111110000000000000000000000000000000000000000000000000000111111111100000000000000000000011111111110000000000000000000000000000001111111111100000000000000001111111111000000000000000000000000000000000000000000000000000011111111110000000000000000000001111111111000000000000000000000000000000111111111110000000000000000111111111100000000000000000000000000000000000000000000000000001111111111000000000000000000000111111111100000000000000000000000000000001111111111000000000000000111111111110000000000000000000000000000000000000000000000000000111111111100000000000000000000011111111100000000000000000000000000000000111111111110000000000000011111111110000000000000000000000000000000000000000000000000000011111111110000000000000000000001111111110000000000000000000000000000000011111111111000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000111111111000000000000000000000000000000001111111111100000000000000111111111100000000000000000000000000000000000000000000000000000111111111100000000000000000000011111111100000000000000000000000000000000111111111110000000000000111111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000001111111100000000000000000000000000000000011111111111100000000000011111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000111111110000000000000000000000000000000001111111111110000000000001111111111100000000000000000000000000000000000000000000000000000011111111000000000000000000000111111111000000000000000000000000000000000111111111111000000000000111111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111100000000000000000000000000000000001111111111100000000000011111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000111111111110000000000001111111111100000000000000000000000000000000000000000000000000000011111111100000000000000000001111111110000000000000000000000000000000000011111111111000000000000111111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111000000000000000000000000000000000001111111111100000000000011111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111100000000000000000000000000000000000011111111110000000000001111111111100000000000000000000000000000000000000000000000000000001111111110000000000000000001111111110000000000000000000000000000000000001111111111100000000000111111111110000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000111111110110000000000011111111111000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000000000000000000000001111111111100000000011111111111000000000000000000000000000000000000000000000000000000001111111110000000000000000111111111100000000000000000000000000000000000000111111111110000000001111111111110000000000000000000000000000000000000000000000000000000111111111100000000000000001111111110000000000000000000000000000000000000001111111111100000000111111111001000000000000000000000000000000000000000000000000000000011111111110000000000000001111111110000000000000000000000000000000000000000111111111110000000011111111101100000000000000000000000000000000000000000000000000000001111111111100000000000001111111111000000000000000000000000000000000000000011111111111000000001111111110110000000000000000000000000000000000000000000000000000000111111111110000000000001111111111100000000000000000000000000000000000000001111111111100000000111111111011000000000000000000000000000000000000000000000000000000011111111111100000000000111111111110000000000000000000000000000000000000000111111111111000000111111111101100000000000000000000000000000000000000000000000000000000111111111110000000000011111111111000000000000000000000000000000000000000011111111111110000011111111110110000000000000000000000000000000000000000000000000000000011111111111000000000011111111111100000000000000000000000000000000000000000111111111111000001111111111011000000000000000000000000000000000000000000000000000000001111111111110000000011111111111100000000000000000000000000000000000000000011111111111110000111111111101100000000000000000000000000000000000000000000000000000000111111111111100000011111111111110000000000000000000000000000000000000000001111111111111000111111111111110000000000000000000000000000000000000000000000000000000011111111111110000011111111111111000000000000000000000000000000000000000000111111111111100011111111111111100000000000000000000000000000000000000000000000000000001111111111111100001111111111111100000000000000000000000000000000000000000011111111111111101111111111111110000000000000000000000000000000000000000000000000000000111111111111110001111111111111110000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111111100111111111111111000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111000111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111000110011111111111000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111110011111111111111100000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111111111111010000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000110000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000011110000001111111111111111111111111111110000000001111111110000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000011011100000111111111111111111111111111111000000111111111111110000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000001000001100011111111111111111111111111111100001111111010111000100000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000001001111111111111111111111111111110001111100000011100000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000110000000110111111111111111111111111111111001110000000001000011100000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000010000000011111111111111111111111111111111101110000000011100001110000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000100000011101111111111111111111111111111110111000000011111101110000000000000000001111000000000000001111111111111111111111111111100000011111100000000000000000000011000110110111111111111111111111111111111111110000011001001000010000000000000001111111110000000000111111111111111111111111111110000111111111000000000000000000101111001001011111111111111111111111111111111111000010000000011111100000000000000111111111100000000011111111111111111111111111111000111111111100000000000000000000111100011101111111111111111111111111111111111000001000000000111110000000000000111111111111100000000111111111111111111111111111100111111111110000000000000000000011010000111111111111111111111111111111111111100001000000000001111000000000000011111111111111000000011111111111111111111111111110011111111111100000000000000000000000000011111111111111111111111111111111111110000100000000000011100000000000011111111111111100000001111111111111111111111111111011111111111000000000000000000000000000011111111111111111111111111111111111111100110000000000000110000000000011000011111111111000001111111111111111111111111111111111111110001100000000000000000000000111111111111111111111111111111111111111110010000000000000000000000000001000000011111111110000111111111111111111111111111111111111111000010000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000011111111110011111111111111111111111111111111111100000001000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000011000000011111111111001111111111111111111111111111111111110001000010000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000011100001111111111111111111111111111111111111111111111111000100001000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000001100111000011111111111111111111111111111111111111111111111000010000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000111100010000111111111111111111111111111111111111111111111100000001110000000000000000000000111111111111111111111111111111111111111110000000000000000000000000000000111101000001111111111111111111111111111111111111111111110000000010000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000010110100000011111111111111111111111111111111111111111110000010101000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000001011010000000111111111111111111111111111111111111111110000001010100000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000101000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000011111111011111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111110011110111011111111111111011111000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000001111111000001001001011111011110000111000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000111111100000000100001111101111000011100000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111100001111001111110111001101100000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000111011111000111111111111111101110110000000000000000000000000000000000000000000000111111111000000111111000000000000000000000000000000000000000000000000000000000001100111110011111111111111101111010000000000000000000000000000000000000000000000001111111111110010110000000000000000000000000000000000000000000000000000000000000010001111111111111111111110111111000000000000000000000000000000000000000000000000000100101111100000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111000000000000000000000000000000000000000000000000000000000101111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000011110010110000000000000000000000000000000000000000000000000000000000000000000000000111111111101111000000000000000000000000000000000000000000000000000000000000000110011100000000000000000000000000000000000000000000000000000000000000000000000000011111110000111100000000000000000000000000000000000000000000000000000000000000000111001000000000000000000000000000000000000000000000000000000000000000000000000001111111111001110000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000100000011100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110011100111000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001100011100000000000000000000000000000000000000000000000000000000000110111110111010000000000000000000000000000000000000000000000000000000000000000000000001111000000001110000000000000000000000000000000000000000000000000000000000011011111011101000000000000000000000000000000000000000000000000000000000000000000000000111001000011111000000000000000000000000000000000000000000000000000000000001110010000111100000000000000000000000000000000000000000000000000000000000000000000000011101111001111000000000000000000000000000000000000000000000000000000000000111110000000010000000000000000000000000000000000000000000000000000000000000000000000001111111110111100000000000000000000000000000000000000000000000000000000000001111100000111000000000000000000000000000000000000000000000000000000000000000000000000111111110000110000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000011111000000111000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000001111110111111100000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end
            STATE_HI2:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_HI1;
						TRANSITION_ME: next_state <= STATE_HI1;
						TRANSITION_HI: next_state <= STATE_HI3;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b100;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000000000000000011111111100000000000000000000001111111100000000000000000000000000000111111111110000000000001111111110000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000111111110000000000000000000000000000011111111111000000000000111111111000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000011111111000000000000000000000000000001111111111100000000000111111111100000000000000000000000000000000000000000000000000000000000011111111100000000000000000000011111111100000000000000000000000000000111111111110000000000011111111110000000000000000000000000000000000000000000000000000000000001111111110000000000000000000001111111110000000000000000000000000000011111111111000000000001111111111000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000111111111000000000000000000000000000001111111111100000000000111111111100000000000000000000000000000000000000000000000000000000000011111111100000000000000000000011111111000000000000000000000000000000011111111110000000000011111111110000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111100000000000000000000000000000001111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000011111111100000000000000000000111111110000000000000000000000000000000011111111111000000000011111111110000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111000000000000000000000000000000001111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111100000000000000000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111110000000000000000000000000000000001111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000111111110000000000000000000111111111000000000000000000000000000000000111111111110000000001111111111000000000000000000000000000000000000000000000000000000000000011111111000000000000000000011111111000000000000000000000000000000000011111111111000000000111111111100000000000000000000000000000000000000000000000000000000000001111111100000000000000000001111111100000000000000000000000000000000001111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000111111110000000000000000000111111110000000000000000000000000000000000111111111110000000001111111111000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111110000000000000000000000000000000000001111111101100000000111111111100000000000000000000000000000000000000000000000000000000000001111111110000000000000000011111111000000000000000000000000000000000000111111110010000000011111111110000000000000000000000000000000000000000000000000000000000000111111111000000000000000011111111100000000000000000000000000000000000011111111101000000001111111111000000000000000000000000000000000000000000000000000000000000011111111100000000000000001111111110000000000000000000000000000000000000111111111100000001111111111100000000000000000000000000000000000000000000000000000000000001111111111000000000000001111111110000000000000000000000000000000000000011111111110000000111111111110000000000000000000000000000000000000000000000000000000000000111111111100000000000000111111111000000000000000000000000000000000000001111111111100000011111111111000000000000000000000000000000000000000000000000000000000000001111111111000000000000111111111100000000000000000000000000000000000000111111110110000001111111111100000000000000000000000000000000000000000000000000000000000000111111111100000000000011111111110000000000000000000000000000000000000011111111001100000111111111110000000000000000000000000000000000000000000000000000000000000011111111110000000000011111111111000000000000000000000000000000000000001111111100110000011111111111000000000000000000000000000000000000000000000000000000000000001111111111100000000001111111111100000000000000000000000000000000000000111111100011000001111111111100000000000000000000000000000000000000000000000000000000000000111111111110000000001111111111110000000000000000000000000000000000000011111110001110000111111111110000000000000000000000000000000000000000000000000000000000000011111111111100000001111111111110000000000000000000000000000000000000001111111001111000111111111111000000000000000000000000000000000000000000000000000000000000001111111111110000001111111111111000000000000000000000000000000000000000111111100111100011111111111100000000000000000000000000000000000000000000000000000000000000111111111111100001111111111111100000000000000000000000000000000000000011111100001110001111111111110000000000000000000000000000000000000000000000000000000000000011111111111110000111111111111110000000000000000000000000000000000000001111111000111101111111111111000000000000000000000000000000000000000000000000000000000000001111111111111000011111111111111000000000000000000000000000000000000000111111100111110111111111111100000000000000000000000000000000000000000000000000000000000000111111111111110011111111111111100000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111100111111111111111000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111100001111111111111000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111100011001111111111000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000111100000000001111111111111111111111111111100000000001111110000000000000000000000000000000000000000000000011111111111111111111111111110000000001111100000000000011111000000000111111111111111111111111111110000000011111111000000000000000000000000000000000000000000000001111111111111111111111111111000000001111110000000000011111000000000011111111111111111111111111111000000111100111110000000000000000000000000000000000000000000000111111111111111111111111111100000001111111100000000001111000001110011111111111111111111111111111100000111100011111000000000000000000000000001111110000000000000011111111111111111111111111100000011111111110000000000111000000111101111111111111111111111111111110111111100000001110000000000000000000000001111111110000000000001111111111111111111111111110000011111111111000000000011100000011111111111111111111111111111111111111111100000000011100000000000000000000000111111111111000000000111111111111111111111111111000111111111111110000000001100000001111111111111111111111111111111111111111110000000000110000000000000000000000011111111111111000000011111111111111111111111111101111111111111111000000000110000001111111111111111111111111111111111111111111100000000000100000000000000000000011111111111111111000011111111111111111111111111111111111111111111100000000010000011111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000001000011111111111111111111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000100000111111111111111111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111011111100000000010000011111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110001111110000000001000000111111111111111111111111111111111111111111111000000000000000000000000000000000111111101111111111111111111111111111111111111111111111111000011111000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000011111100011111111111111111111111111111111111111111111110000001111100000000000000000111111111111111111111111111111111111111111000000000001111100000000000000000001111110000011111111111111011110111111111111111111111111000000111100000000000000000001111111111111111111111111111111111111111100000000000011110000000000000000000111111000000011111111110001111011011111111111110011111100000011110000000000001000000011111111111111111111111111111111111111100000000000001110000000000000000000001111100000000111111111000000000100101111011111001111100000001111000000000001110000000111111111111111111111111111111111111100000000000001100000000000000000000000111110000000001111111010000000010000111101110000111100000000111100000000000111000000001111111111111111111111111111111111100000000000001000000000000000000000000011111000000000011111100000000011001111110011000001110000000110000000000000100110000000011111111111111111111111111111111100000000000000000000000000000000000000001111100000000000111110011000011111111111000000000110000000100000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000011000000000000111000000011111111111110000010010000000000000000000000000000000000000000001111111111000011111111110000000000000001000000000000000000000000000000000010000000000001100111101111111111111001111000000000000000000000000000000000010000000000001111111111100111100000000000000000000000000000000000000000000000000000000000000000000010111111111111111111111110000000000100000000000000000000000000000000000000001001011110001100000000000000000000000000010100000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000101000000000000000000000000011111100000000000000000000000000000101010000000000000000000000000000100000000000000000011111111111111100000000000000000000000000000010101000000000000000000000001111111000000000000000000000000001010101000000000000000000000000000000000000000000000000111111111111110000000000000000000010100000001010100100000000000000000001111111100000000000000000000000000001010000000000000000000000000000000000000000000000000001111111111111000000000000000000101010000000001010000000000000000000000111111111000000000000000000000000000101000000000000000000000000000000000000000000000000000111100000111100000000000000010010101000000000101000000000000000000000001100100010000000000000000000000000010000000000000000000000101000000000000000000000000000011111110011110000000000000000001010100000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000010101000000000000000000000000001111110001111000000000000000000101000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000001010100100000000000000000000000111111111111100000000000000000010100000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000001010000000000000000000000000011110110001111000000000000000001000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000101000000000000000000000000001100011100011100000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000011110000000000000000000000000000000000000000000000000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000111111000000000000000000000000000000000000000000000000000000110111100111000000000000000000000000000000000000000000000000000000000000000000000000000000011011110111111000000000000000000000000000000000000000000000000000000011001110011101000000000000000000000000000000000000000000000000000000000000000000000000000000111111011111100000000000000000000000000000000000000000000000000000001110000000010100000000000000000000000000000000000000000000000000000000000000000000000000000111111000001110000000000000000000000000000000000000000000000000000000011110000000110000000000000000000000000000000000000000000000000000000000000000000000000000001110000001111000000000000000000000000000000000000000000000000000000001111100011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100100111000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end
            STATE_HI3:begin
                    case (transition)
						TRANSITION_LO: next_state <= STATE_HI2;
						TRANSITION_ME: next_state <= STATE_HI2;
						TRANSITION_HI: next_state <= STATE_HI2;
						default: next_state <= current_state;
					endcase
					color_background_reg <= 3'b100;
					color_foreground_reg <= 3'b111;
					current_image <= 19200'b000000000000000000000000000000000000000111111110000000000111111110000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000011111111000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000001111111110000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111000000000000000000000000000000111111111100000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111100000000000000000000000000000011111111110000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110000000000000000000000000000001111111111000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000011111111000000000000000000000000000000111111111100000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000001111111000000000000000000000000000000011111111110000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000111111100000000000000000000000000000001111111111000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000011111110000000000000000000000000000000111111111100000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000011111111000000000000000000000000000000011111111110000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000001111111100000000000000000000000000000001111111111000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111110000000000000000000000000000000111111111100000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000011111110000000000000000000000000000000001110111110000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000001111111000000000000000000000000000000000111111111100000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000111111100000000000000000000000000000000011111110110000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000000000000000000000000001111111111000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000011111111000000000000000000000000000000000111111111100000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000001111111100000000000000000000000000000000011111111111000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000001111111110000000000000000000000000000000001111111111100001111111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000111111111000000000000000000000000000000000111111111111000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111100000000000000000000000000000000001111111111100111111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000011111111110000000000000000000000000000000000111111111110011111111110100000000000000000000000000000000000000000000000000000000000000000000000000001111111111000011111111111000000000000000000000000000000000011111111111001111111111010000000000000000000000000000000000000000000000000000000000000000000000000000111111111110001111111111100000000000000000000000000000000001111111111110111111111101000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000111111111110000000000000000000000000000000000111111111111011111111110100000000000000000000000000000000000000000000000000000000000000000000000000011111111111100111111111111000000000000000000000000000000000011111111111101111111111010000000000000000000000000000000000000000000000000000000000000000000000000001111111111111011111111111100000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111101111111111110000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111111111111000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111000111111111111000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111000100011111111100000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111111111110000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000001111111111111111110111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111100111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000011100011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111000000111000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000010000001111111111111111111111111111111111111111111100000001100000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111111111011111111111111111111111110000000000000000111111111111111111111111111111111111111111111100010000000000000000000000000000000000000000000000000111111111111111111100011101111111111111111111110000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000001111111111111111001110001010101111111111111111111100000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111111111000000100101011111111111111111111111100000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111110000011110111111110111111111111111111000000000000000011111111111111000111111111111111000000000000000000000000000000000000000000000000000000111111111111111111110001101111111111111001111111111111111110000000000000000000000011110000000110000000000000000000000000000000000000000000000000000000000000000111111111111111111111001111111111111111100111111111111111111000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111101111111111111111100010000000111111111100000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000011111111111100000000000000111111110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000001111111111100000000000000001111111000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000111111111110000000000000000111111100000000000000000000000000111001101000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000011100001111000000000000000011111110000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001110110011100000000000000001111110000000000000000000000000000001100100000000000000000000000001100000000000000000000000000000000000000111111100000000000000000000111111001111000000000000000111111000000000000000000000000000000001000000000000000000000000000101100000000000000000000000000000000000011111110000000000000000000111100001111100000000000000011111100000000000000000000000001100000100000000000000000000000000000010000000000000000000000000000000000001111111000000000000000000011001110001110000000000000001111110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000001100000000111000000000000001111111000000000100000000000000011001110111000000000000000000000000000000000000000000000000000000000000000001111110000000000000000001111100001111100000000000000111111000000000000000000000000001110111011000000000000000000000100011000000000000000000000000000000000000000111111000000000000000000111111011111110000000000000011111001010001000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000011111101111110000000000000001111100001010100000000000000000001111000000110000000000000000000000000000000000000000000000000000000000000001111110000000000000000000110000000111000000000000000100100000001010000000000000000000111110001111000000000000000000000101010000000000000000000000000000000000000110000000000000000000000011100000111000000000000000110000000000100000000000000000000001111111111100000000000000000001010101000000000000000000000000000000000000011000000000000000000000001111111111100000000000000010000000000010000000000000000000000011111111110000000000000000000101010000000000000000000000000000000000000000000000000000000000000000011111111100000000000000001000000000000000000000000000000000000011111111000000000000000000010100000000000000000000000000000000000000000000000100000000000000000001111111100000000000000001100000000000000000000000000000000000000011110000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000011111110000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000111000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                end
            default: next_state = current_state;
        endcase
    end // state_table
    
    // State Registers
    always @(posedge CLOCK_50)
    begin
        if(resetn == 1'b0)
            current_state <= INITIAL_STATE;
        else
            current_state <= next_state;
    end

	wire [2:0] color;
	wire [7:0] x;
	wire [6:0] y;

	reg on_reg;

	always @(posedge CLOCK_50)
		on_reg <= 1'b1;

	wire on;
	assign on = on_reg;

	vga_adapter VGA(
		.resetn(resetn),
		.clock(CLOCK_50),
		.colour(color),
		.x(x),
		.y(y),
		.plot(on),
		/* Signals for the DAC to drive the monitor. */
		.VGA_R(VGA_R),
		.VGA_G(VGA_G),
		.VGA_B(VGA_B),
		.VGA_HS(VGA_HS),
		.VGA_VS(VGA_VS),
		.VGA_BLANK(VGA_BLANK_N),
		.VGA_SYNC(VGA_SYNC_N),
		.VGA_CLK(VGA_CLK)
	);
	defparam VGA.RESOLUTION = "160x120";
	defparam VGA.MONOCHROME = "FALSE";
	defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
	defparam VGA.BACKGROUND_IMAGE = "black.mif";

	imageprocessor ip(
		// Input
		.clock(CLOCK_50),
		.resetn(resetn),
		.image(image),
		.color_background(color_background),
		.color_foreground(color_foreground),
		// Output
		.x(x),
		.y(y),
		.color(color)
	);

    // Debugging Output
    assign LEDR[3:0] = current_state;
	assign LEDG[1:0] = transition;
	segment_decoder seg0(.c(buff[3:0]), .h(HEX0));
	segment_decoder seg1(.c(buff[7:4]), .h(HEX1));
	segment_decoder seg2(.c(buff[11:8]), .h(HEX2));
	segment_decoder seg3(.c(buff[15:12]), .h(HEX3));
	segment_decoder seg4(.c(buff[19:16]), .h(HEX4));
	segment_decoder seg5(.c(buff[23:20]), .h(HEX5));
	segment_decoder seg6(.c(buff[27:24]), .h(HEX6));
	segment_decoder seg7(.c(buff[31:28]), .h(HEX7));
endmodule

